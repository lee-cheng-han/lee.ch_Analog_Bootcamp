** sch_path: /home/leech/lee.ch_Analog_Bootcamp/analog/schematics/testbenches/tb_outimpedence.sch
**.subckt tb_outimpedence VOUT
*.opin VOUT
x1 net1 VOUT net3 GND net2 opamp_single_stage
VDD net1 GND 1.8
VSS net2 GND 0
V1 net3 GND dc 0.9 ac 0
I0 GND VOUT dc 0 ac 1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/leech/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/leech/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/leech/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/leech/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.ac dec 10 1 10G
.control
run
let zout = abs(v(vout))
meas ac Zout_cl MAX zout FROM=1 TO=10
.endc




**** end user architecture code
**.ends

* expanding   symbol:  opamp_single_stage.sym # of pins=5
** sym_path: /home/leech/lee.ch_Analog_Bootcamp/analog/schematics/opamp_single_stage.sym
** sch_path: /home/leech/lee.ch_Analog_Bootcamp/analog/schematics/opamp_single_stage.sch
.subckt opamp_single_stage VDD VOUT VIN_P VIN_N VSS
*.ipin VDD
*.ipin VIN_P
*.ipin VSS
*.opin VOUT
*.ipin VIN_N
XM4 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 VIN_N net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 VIN_P net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VOUT net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 net5 VOUT sky130_fd_pr__cap_mim_m3_1 W=25 L=20 MF=1 m=1
XM8 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1.0 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net3 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1.0 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 VOUT net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1.0 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 net5 net2 7k m=1
XR2 net4 VDD VDD sky130_fd_pr__res_high_po W=0.35 L=14 mult=1 m=1
.ends

.GLOBAL GND
.end
